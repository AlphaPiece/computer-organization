//SW[2:0] data inputs
//SW[9] select signal
//LEDR[0] output display

module mux2to1(SW, LEDR);
    input [9:0] SW;
    output [9:0] LEDR;

    mux_2_1 u0(
        .x(SW[0]),
        .y(SW[1]),
        .s(SW[9]),
        .m(LEDR[0])
        );

endmodule

module mux_2_1(x, y, s, m);
    input x; //selected when s is 0
    input y; //selected when s is 1
    input s; //select signal
    output m; //output
  
    assign m = s & y | ~s & x;
    // OR
    // assign m = s ? y : x;

endmodule
